-- Exercise 3.27
-- logic function

library ieee;
use ieee.std_logic_1164.all;

entity foo is
  port(x, y, z : in std_logic; 
       output : out std_logic);
end foo;

architecture impl of foo is
begin


   -- Add your code here (start)
   output <= ...;
   -- Add your code here (end)
   
   
   
end impl;